module halfAdder (a, b, s, c);
    
    input a, b;
    output logic s, c;

    always_comb begin: 
        s = a ^ b;
        c = a & b;
    end

endmodule: halfAdder

